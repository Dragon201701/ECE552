module pipeline (flush, stall);
	output flush, stall;
	assign flush = 1'b0;
	assign stall = 1'b0;
endmodule