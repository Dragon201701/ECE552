module mux8_16 ();
	input	[2:0]	sel;
	input	[15:0]	in0, in1, in2, in3, in4, in5, in6, in7;
	output	[15:0]	out;

endmodule
